library ieee;
use ieee.std_logic_1164.all;

package mytypes is
	
	subtype led_data is std_logic_vector(23 downto 0);
	
end package;

package body mytypes is

end package body;